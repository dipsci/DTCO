// auto build by GRO compiler 09/12/2022 14:04:48
`define DL_NUM       6 // GRO : delay line number
`define SEL_BITS     3 // GRO : select bitwidth
`define RPC_BITS    16 // GRO : ripple counter bitWidth
`define RO_ACTIVE            1 // SPI : ro active flag
`define SPI_CYCLE        3333.3 // SPI : controller clock period
`define SPI_DWIDTH          16 // SPI : bitWidth
`define INT_CYCLE        1000.0 // SPI : internal clock period
`define PAT_NUM             10 // SPI : number of patterns
`define GRO_CYCLE         10.0 // SPI : GRO clock period
`define RO_GRID_NUM         16 // SPI : number of ro
`define RO_EN_COUNT_BITS     8 // SPI : ro enable count bitwidth
